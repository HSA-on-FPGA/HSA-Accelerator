--
-- Copyright 2017 Konrad Haeublein
--
-- konrad.haeublein@fau.de
--
-- This program is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.
--



-- Content: Kernel File
-- OP-ID : 0
-- This file has been generated by pipegen
-- www3.cs.fau.de
-- konrad.haeublein@fau.de
-- Creation Date: 2017-01-19T12:40:01.697+01:00

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.pkg_custom_config.all;

entity op_0_kernel is
generic(
  g_ivaluewidth : natural:= c_ival_op_0;
  g_ovaluewidth : natural:= c_oval_op_0;
  
  g_windowwidth : natural:= c_ww_op_0;
  g_windowheight: natural:= c_wh_op_0;
  
  g_dummy : natural:= 0
);
port(
  clk   : in std_logic;
  rst_n : in std_logic;
  en    : in std_logic;
  nd    : in std_logic;
  
  di0   : in  std_logic_vector(g_windowwidth*g_windowheight*g_ivaluewidth-1 downto 0);
    
  do0 : out  std_logic_vector(g_ovaluewidth-1 downto 0);
  
  
  valid : out std_logic 
);
end op_0_kernel;

architecture behavior of op_0_kernel is


type VEC_DIN is array (0 to g_windowwidth*g_windowheight-1) of std_logic_vector(g_ivaluewidth-1 downto 0);
signal s_di : VEC_DIN;
signal s_read : std_logic_vector(g_windowwidth*g_windowheight-1 downto 0); 
  
signal s_do_write : std_logic_vector(1-1 downto 0);
signal s_empty_n, s_start, s_do_full, s_done, s_idle, s_rst, s_ready : std_logic;

begin

sig_gen: for i in 0 to g_windowwidth*g_windowheight-1 generate
	s_di(i) <= di0((i+1)*g_ivaluewidth-1 downto i*g_ivaluewidth);
end generate;

s_start <= nd and en;
s_rst <= not rst_n;

process(s_start)
begin
  if s_start='1' then
    s_empty_n <= '1';
    s_do_full <= '1';
  else
    s_empty_n <= '0';
    s_do_full <= '0';
  end if;
end process;

hls_kernel: entity work.kuwahara
port map (
 
  din0_0_V => s_di(0),

       
  din0_1_V => s_di(1),

       
  din0_2_V => s_di(2),

       
  din0_3_V => s_di(3),

       
  din0_4_V => s_di(4),

       
  din0_5_V => s_di(5),

       
  din0_6_V => s_di(6),

       
  din0_7_V => s_di(7),

       
  din0_8_V => s_di(8),

       
  din0_9_V => s_di(9),

       
  din0_10_V => s_di(10),

       
  din0_11_V => s_di(11),

       
  din0_12_V => s_di(12),

       
  din0_13_V => s_di(13),

       
  din0_14_V => s_di(14),

       
  din0_15_V => s_di(15),

       
  din0_16_V => s_di(16),

       
  din0_17_V => s_di(17),

       
  din0_18_V => s_di(18),

       
  din0_19_V => s_di(19),

       
  din0_20_V => s_di(20),

       
  din0_21_V => s_di(21),

       
  din0_22_V => s_di(22),

       
  din0_23_V => s_di(23),

       
  din0_24_V => s_di(24),

       
  ap_return => do0,

  ap_clk  => clk,
  ap_rst  => s_rst,
  ap_done => s_done,
  ap_start => s_start,
  ap_idle => s_idle,  
  ap_ready => s_ready
);
     
valid <= s_done;

end behavior;

     
