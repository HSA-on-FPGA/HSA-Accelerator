--
-- Copyright 2017 Konrad Haeublein
--
-- konrad.haeublein@fau.de
--
-- This program is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.
--

-- Content: Config File
-- This file has been generated by pipegen
-- www3.cs.fau.de
-- konrad.haeublein@fau.de
-- Creation Date: 2017-01-19T12:40:00.973+01:00


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.pkg_config.all;

package pkg_custom_config is
---------------------------------------
------- Generated Parameters ----------
---------------------------------------
constant c_picwidth  : integer:= 128;
constant c_picheight : integer:= 128;
constant c_ctrlwidth : integer:= 1;  

---- Kernel Parameters ---


--- Constant Definition of Kernel_0 ---


-- only width of buffer gray supported
constant c_ival_op_0 : integer:= c_dw_pix_max_gray_0; 
constant c_oval_op_0 : integer:= c_dw_pix_max_gray_0; -- Must be equal to ival in case c_ic > 1

constant c_ww_op_0 : integer:= c_ww_max_0;  
constant c_wh_op_0 : integer:= c_wh_max_0;   
constant c_kd_op_0: integer:= 1; -- Kernel delay for defining ctrl channel, not relevant
constant c_ic_op_0 : integer:= 1; -- Number of kernel iterations

---------------------------------------------
-------- End of Generated Parameters --------
---------------------------------------------

--- Required for Testbench ---
constant picsize : integer:= c_picwidth*c_picheight;


end pkg_custom_config;

