--
-- Copyright 2017 Konrad Haeublein
--
-- konrad.haeublein@fau.de
--
-- This program is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.pkg_functions.all;

package pkg_config is
--------------------------------------------
------- Parameters for Accelerator_PE_0 ----
--------------------------------------------

-- Global Configurable Parameters --

--- Values for maximum config settings and structural parameters

-- Following Value can have artibrary confifugration

constant c_iw_max_0   : integer:= 4100; -- Maximum image width
constant c_ih_max_0   : integer:= 4100; -- Maximum image height

constant c_ww_max_0   : integer:= 5; -- Maximum window width
constant c_wh_max_0   : integer:= 5; -- Maximum window height

constant c_ww_min_0   : integer:= 2; -- Minimum window width
constant c_wh_min_0   : integer:= 2; -- Minimum window height

constant c_dw_pix_max_0   : integer:= 8; -- Maximum datawith for pixel in RGB channel, should be 8 for current tb
constant c_dw_pix_max_gray_0 : integer:= 16; -- Maximum datawith for pixel in gray channel, must be equal or higher than pix_max!
constant c_num_col_max_0 : integer:= 3; -- Maximum number of supported colors, should be 3 for current tb

constant c_par_0  : integer:= 1  ; -- Factor for Vectorization! 
constant c_en_border_handling_0 : boolean:= true; -- if true bits for border handling are respected
constant c_num_custom_kernel_0 : integer:= 0; -- if 1, custom kernel, generated by vivado HLS will be used

---------------------------------------------------------------------
-- ALL Following Values may NOT be changed for current AXI wrapper!!!!
---------------------------------------------------------------------

-- Structural Parameters

constant c_it_0  : integer:= 1; -- should be changed at one time
constant c_num_kernel_0 : integer:= 3; -- Total number of Kernel modules
constant c_num_kmodes_0 : integer:= 5; -- Total number of supported operations
constant c_num_bmodes_0 : integer:= 3; -- Total number of supported  border handling operations
constant c_num_im_para_0 : integer:= 8; -- Total number of image parameters



--------------------------------------------------------------

----             Operation Register: Addr=5
--               ------------------------------------------------------
--   Descripiton | Reserved|Color|   Border   |   Kernel   |Norm/Tresh|
--               ------------------------------------------------------

--  Num of Bits      ...   |  1  |     2      |        3   |     1    |
--  Decoding    --------------------------------------------------------
--     0                   |Color|     Off    |Single Conv.|   Off    |
--     1                   |Gray |   Zero Pad |Dual Conv.  |   On     |
--     2                   |     |   Clamp    |Median      |          |
--     3                   |     |            |Erosion     |          |
--     4                   |     |            |Dilation    |          |


--- Coding internal Register


-- Register Configuration | Register
------------------------------------
-- Resolution X Dimension  |   0
-- Resolution Y Dimension  |   1
-- Number of Pixel in Image|   2
-- Windowwidth X Dimension |   3
-- Windowwidth Y Dimension |   4
-- Operation               |   5
-- Normalize Value         |   6
-- Treshold Value          |   7
-- Coefficient Value_0     |   8
--            ....         |   ..
-- Coefficient Value_49    |   57

---------------------
--Axi PE_0 ---
----------------------

constant c_numpix_addr_0: integer:= 2; -- address for Number of Pixel Register
constant c_op_addr_0: integer:= 5; -- address for operation
constant c_pack_size_0: integer:= 32; -- counter for TLAST signal in AXI Stream Master
-- constant c_dev_ultra_0: boolean:= false; -- selects fifo xilinx fifo macro for correct device
constant c_rst_interval_0: integer:= 10; -- duration for holding reset 

---------------------
--Accelerator_PE_0 ---
----------------------

constant c_np_max_0 : integer:= c_iw_max_0*c_ih_max_0; -- max number of total pixels
constant c_np_addr_0 : integer:= f_log2(c_np_max_0);

constant c_num_col_chan_0 : integer:= c_num_col_max_0-1;
-- Definition of datawidth, lower values gray uper values other colors (RGB=8+8+16=32)
constant c_dw_pe_0 : integer:= c_num_col_chan_0 * c_dw_pix_max_0 + c_dw_pix_max_gray_0;
-- Total number  of Registers: 7 + 2*5*5;
constant c_num_reg_0 : integer:= c_num_im_para_0 + 2*c_ww_max_0*c_wh_max_0;
constant c_reg_addr_0 : integer:= f_log2(c_num_reg_0);

--type VEC_REG_0 is array(0 to c_num_reg_0-1) of std_logic_vector(c_regw_0-1 downto 0);
type VEC_DCOL_0 is array(0 to c_num_col_chan_0-1) of std_logic_vector(c_par_0*c_dw_pix_max_0-1 downto 0);

type VEC_DPEPAR_0 is array(0 to c_par_0-1) of std_logic_vector(c_dw_pe_0-1 downto 0);

type BORDER_STATE_0 is (up_left, up, up_right, left, right, down_left, down, down_right, no_border);
----------------------
---- Buffer_CLB_0 ----
----------------------

constant c_iw_addr_0 : integer:= f_log2(c_iw_max_0);
constant c_ih_addr_0 : integer:= f_log2(c_ih_max_0);


constant c_ww_addr_0 : integer:= f_log2(c_ww_max_0);
constant c_wh_addr_0 : integer:= f_log2(c_wh_max_0);

type VEC_MASK_0 is array(0 to c_ww_max_0-1) of std_logic_vector(c_dw_pix_max_0-1 downto 0);
type ARRAY_MASK_0 is array(0 to c_wh_max_0-1) of VEC_MASK_0;
type ARRAY_MASKPAR_0 is array(0 to c_par_0-1) of ARRAY_MASK_0;
type ARRAY_MASKPARCOL_0 is array(0 to c_num_col_max_0-1) of ARRAY_MASKPAR_0;


----------------------
---- Buffer_CLB_Gray_0 
----------------------

type VEC_MASK_GRAY_0 is array(0 to c_ww_max_0-1) of std_logic_vector(c_dw_pix_max_gray_0-1 downto 0);
type ARRAY_MASK_GRAY_0 is array(0 to c_wh_max_0-1) of VEC_MASK_GRAY_0;
type ARRAY_MASKPAR_GRAY_0 is array(0 to c_par_0-1) of ARRAY_MASK_GRAY_0;

----------------------
---- Kernel_CLB_0 ----
----------------------

constant c_normw_0 : integer:= c_dw_pix_max_0;
constant c_treshw_0 : integer:= c_dw_pix_max_gray_0;

constant c_kinstrw_0 : integer:= f_log2(c_num_kmodes_0)+1;
constant c_dw_addr_0 : integer:= f_log2(c_dw_pix_max_0);
constant c_coeffw_0 : integer:= c_dw_pix_max_0+1; -- for calulating with signed values

type VEC_KERNEL_0 is array(0 to c_ww_max_0*c_wh_max_0-1) of std_logic_vector(c_dw_pix_max_0-1 downto 0);
type VEC_COEFF_0 is array(0 to c_ww_max_0*c_wh_max_0-1) of std_logic_vector(c_coeffw_0-1 downto 0);


----------------------
---- Kernel_CLB_Gray_0 ----
----------------------

constant c_normw_gray_0 : integer:= c_dw_pix_max_0;
constant c_treshw_gray_0 : integer:= c_dw_pix_max_gray_0;

type VEC_KERNEL_GRAY_0 is array(0 to c_ww_max_0*c_wh_max_0-1) of std_logic_vector(c_dw_pix_max_gray_0-1 downto 0);




end pkg_config;
